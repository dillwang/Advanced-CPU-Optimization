module map_table(
    input clk,
    input rst_n,
    input rename_valid,
    input 
)