module ghr(

input clk,
input rst_n,
input logic branch_outcome,
